module ReservationStation(
   
);

    
    

endmodule