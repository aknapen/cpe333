module ReorderBuffer(
   
);

    
    

endmodule