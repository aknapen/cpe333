module TaskGeneration(
   
);

    
    

endmodule